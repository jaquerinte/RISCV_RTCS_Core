//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define SIM 1

`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Generate random number
// Description  : Generate a random number and send by the output

//***Headers***
`include "defines.vh"
//***Module***
module random_number_generator #(
        parameter integer WORD_SIZE = 32
    )
    (
        input  clk_i ,
        output [WORD_SIZE - 1 : 0] output_number_o 
    );

//***Interal logic generated by compiler***  


//***Dumped Internal logic***
    assign output_number_o =  32'b00000001010000100100101111001001;
    //assign output_number_o = 32'b00100110011111101110111100010000  ;
    
//***Handcrafted Internal logic*** 
//TODO
endmodule

`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Memory emulator for the processor
// Description  : Memory simulation using a 32 bit size and a LINE_SIZE of 128 with a delay in 3 cycles for geting the data
// Coder        : Jaquer AND VORIXO

//***Headers***
`include "defines.vh"
//***Module***
module memory #(
        parameter integer WORD_SIZE = 32,
        parameter integer WORDS_PER_LINES = 4,
        parameter integer LINE_SIZE = 128,
        parameter integer MEMORY_LINES = 32
    )
    (
        input  clk_i ,
        input  rstn_i ,
        input  we_i ,
        input  strobe_i ,
        input  [LINE_SIZE - 1 : 0] data_i ,
        input  [WORD_SIZE - 1 : 0] addr_i ,
        output [LINE_SIZE - 1 : 0] data_o ,
        output valid_data_o 
    );

//***Interal logic generated by compiler***  


//***Dumped Internal logic***
    reg [WORD_SIZE-1:0] main_mem [0:MEMORY_LINES-1];
    reg [LINE_SIZE-1:0] data_o_0;
    reg [LINE_SIZE-1:0] data_o_1;
    reg [LINE_SIZE-1:0] data_o_2;
    reg [LINE_SIZE-1:0] data_o_3; 
    reg [LINE_SIZE-1:0] data_o_4;    
    reg valid_0; 
    reg valid_1;
    reg valid_2;
    reg valid_3;
    reg valid_4;
    `ifdef SIM
        initial begin
        $display("Loading rom.");
        $readmemh("../../../memory.hex", main_mem);
        $display("Rom loaded");
        end
    `endif

    always @(posedge clk_i) begin
        // data_o_0 <= {WORD_SIZE{1'b0}};
        valid_0 <=0;                           
        if (!rstn_i) begin                                       
            // reset                                            
            integer i;         
            /* verilator lint_off BLKLOOPINIT*/                                 
            for(i=0;i<MEMORY_LINES; i=i+1) begin                 
                main_mem[i] <= {WORD_SIZE{1'b0}};                
            end   
            /* verilator lint_on BLKLOOPINIT*/                                             
                                                                
        end                                                  
        else if (we_i) begin                                 
            main_mem[addr_i] <= data_i[31:0] ;                         
                                                                
        end else if (strobe_i) begin                        
            data_o_0[31:0] <=  main_mem[addr_i>>5]; 
            data_o_0[63:32] <= main_mem[(addr_i>>5)+1];
            data_o_0[95:64] <= main_mem[(addr_i>>5)+2];          
            data_o_0[127:96] <= main_mem[(addr_i>>5)+3]; 
            //data_o_0[31:0] <=  main_mem[addr_i];           
            //data_o_0[63:32] <= main_mem[addr_i + 2'b01];
            //data_o_0[95:64] <= main_mem[addr_i + 2'b10];                 
            //data_o_0[127:96] <= main_mem[addr_i + 2'b11]; 
            valid_0 <= 1;                    
                                                                
        end
        data_o <= data_o_4;
        valid_data_o <= valid_4;
        data_o_4 <=  data_o_3;
        valid_4 <= valid_3;
        data_o_3 <= data_o_2;
        valid_3 <= valid_2;
        data_o_2 <= data_o_1;
        valid_2 <= valid_1;
        data_o_1 <= data_o_0;
        valid_1 <= valid_0;

    end   
    
//***Handcrafted Internal logic*** 
//TODO
endmodule

`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND Barrera

//***Headers***
`include "defines.vh"
//***Module***
module processor #(
        parameter integer WORD_SIZE = 32,
        parameter integer REGISTERS = 32,
        parameter integer LINE_SIZE = 128,
        parameter integer ALUOP_SIZE = 4,
        parameter integer REGDIRSIZE = 5
    )
    (
        input  clk_i ,
        input  rstn_i 
    );

//***Interal logic generated by compiler***  
    wire [WORD_SIZE - 1 : 0] addr_IF_MEM; // wiring between addr_o of module IF and addr_i of module MEM
    wire valid_data_MEM_IF; // wiring between valid_data_o of module MEM and valid_input_i of module IF
//***Auxiliar Wires***  
    wire [LINE_SIZE - 1 : 0] mem_data_bus_w; // Auxiliar Wire
    wire write_data_bus_mem_w; // Auxiliar Wire
    wire strobe_main_memory_w; // Auxiliar Wire

    fetch #(
        .WORD_SIZE (32),
        .LINE_SIZE (128),
        .WORDS_PER_LINES (4),
        .MEMORY_LINES (4),
        .TAG (24),
        .OFFSET (7)
    )
    inst_IF(
        .clk_i                        (clk_i ),
        .rstn_i                       (rstn_i ),
        .data_i                       (mem_data_bus_w),
        .valid_input_i                (valid_data_MEM_IF),
        .nrm0_o                       (),
        .addr_o                       (addr_IF_MEM),
        .instruction_register_o       (),
        .ask_memory_o                 (strobe_main_memory_w),
        .valid_o                      ()
    );

    memory #(
        .WORD_SIZE (32),
        .WORDS_PER_LINES (4),
        .LINE_SIZE (128),
        .MEMORY_LINES (32)
    )
    inst_MEM(
        .clk_i                (clk_i ),
        .rstn_i               (rstn_i ),
        .we_i                 (write_data_bus_mem_w),
        .strobe_i             (strobe_main_memory_w),
        .data_i               (mem_data_bus_w),
        .addr_i               (addr_IF_MEM),
        .data_o               (mem_data_bus_w),
        .valid_data_o         (valid_data_MEM_IF)
    );


//***Handcrafted Internal logic*** 
//TODO
endmodule

`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Generate the hash function
// Description  : Generate all function

//***Headers***
`include "defines.vh"
//***Module***
module hash_cache_function #(
        parameter integer WORD_SIZE = 32
    )
    (
        input  clk_i ,
        input  [WORD_SIZE - 1 : 0] addr_i ,
        output line_index_o 
    );

//***Interal logic generated by compiler***  
//***Auxiliar Wires***  
    wire [WORD_SIZE - 1 : 0] random_number_w; // Auxiliar Wire

    random_number_generator #(
        .WORD_SIZE (32)
    )
    inst_RNG(
        .clk_i                  (clk_i ),
        .output_number_o        (random_number_w)
    );


//***Dumped Internal logic***
    reg [WORD_SIZE-1:0] rotate_0;
    reg [WORD_SIZE-1:0] rotate_1;
    reg [WORD_SIZE-1:0] rotate_2;
    reg [WORD_SIZE-1:0] rotate_3;
    reg [WORD_SIZE-1:0] rotate_4;
    reg [WORD_SIZE-1:0] rotate_5;
    wire [(WORD_SIZE*3)-1:0] output_xor_0;
    wire [48-1:0] output_xor_1;
    wire [24-1:0] output_xor_2;
    wire [12-1:0] output_xor_3;
    wire [6-1:0] output_xor_4;
    wire [3-1:0] output_xor_5;
    wire output_xor_6;
    

    assign output_xor_0 = {rotate_0,rotate_1,rotate_2} ^ {rotate_3,rotate_4,rotate_5};
    assign output_xor_1 = output_xor_0[95:48] ^ output_xor_0[47:0];
    assign output_xor_2 = output_xor_1[47:24] ^ output_xor_1[23:0];
    assign output_xor_3 = output_xor_2[23:12] ^ output_xor_2[11:0];
    assign output_xor_4 = output_xor_3[11:6] ^ output_xor_3[5:0];
    assign output_xor_5 = output_xor_4[5:3] ^ output_xor_4[2:0];
    assign line_index_o = output_xor_5[2] ^ output_xor_5[1] ^ output_xor_5[0];

    always @(posedge clk_i) begin


    rotate_0  <= (random_number_w >> addr_i[11:7]) | (random_number_w <<  (WORD_SIZE - {{27{1'b0}},addr_i[11:7]}));
    rotate_1  <= (random_number_w >> addr_i[16:12]) | (random_number_w <<  (WORD_SIZE - {{27{1'b0}},addr_i[16:12]}));
    rotate_2  <= (random_number_w >> addr_i[21:17]) | (random_number_w <<  (WORD_SIZE - {{27{1'b0}},addr_i[21:17]}));

    rotate_3  <= ({addr_i[31:7],7'b0000000} >> random_number_w[4:0]) | ({addr_i[31:7],7'b0000000} <<  (WORD_SIZE - {{27{1'b0}},random_number_w[4:0]}));
    rotate_4  <= ({addr_i[31:7],7'b0000000} >> random_number_w[9:5]) | ({addr_i[31:7],7'b0000000} <<  (WORD_SIZE - {{27{1'b0}},random_number_w[9:5]}));
    rotate_5  <= ({addr_i[31:7],7'b0000000} >> random_number_w[14:10]) | ({addr_i[31:7],7'b0000000} <<  (WORD_SIZE - {{27{1'b0}},random_number_w[14:10]}));



    end


    
//***Handcrafted Internal logic*** 
//TODO
endmodule
